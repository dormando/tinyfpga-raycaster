// (modified heavily) from mojo example source code.
// (same MIT license)

// NOTE: original module didn't work with CLK_DIV=1 (half clock)
// I've cut out a bunch of it, breaking MOSI.
// it's fixable but I'm not currently using it.
// CPOL/CPHA 0

module spi #(parameter CLK_DIV = 2)(
    input clk,
    input rst,
    input miso,
    output reg mosi,
    output reg sck,
    input start,
    output reg ss, // lcd_ss
    input[7:0] data_in,
    output[7:0] data_out,
    output busy,
    output new_data
);

localparam STATE_SIZE = 2;
localparam IDLE = 2'd0,
           WAIT_HALF = 2'd1,
           TRANSFER = 2'd2;

reg [STATE_SIZE-1:0] state_d, state_q;

reg [7:0] data_d, data_q;
reg sck_d, sck_q;
reg mosi_d, mosi_q;
reg [2:0] ctr_d, ctr_q;
reg new_data_d, new_data_q;
reg [7:0] data_out_d, data_out_q;

assign busy = state_q != IDLE;
assign data_out = data_out_q;
assign new_data = new_data_q;

always @(*) begin
    data_d = data_q;
    ctr_d = ctr_q;
	new_data_d = 1'b0;
	data_out_d = data_out_q;
	state_d = state_q;
    ss = 1'b0; // ss low when active.
    sck = 1'b0;
    mosi = 1'b0;

    case (state_q)
        IDLE: begin
            sck_d = 4'b0;
            ctr_d = 3'b111;
            ss = 1'b1; // high when idle.
            if (start == 1'b1) begin
                data_d = data_in;
                state_d = WAIT_HALF;
            end
        end
        WAIT_HALF: begin
            sck = 1'b0;
            mosi = data_q[ctr_q];
            state_d = TRANSFER;
        end
        TRANSFER: begin
            sck = 1'b1;
            mosi = data_q[ctr_q];
            ctr_d = ctr_q - 1'b1;
            if (ctr_q == 3'b000) begin
                state_d = IDLE;
                data_out_d = data_q;
                new_data_d = 1'b1;
            end else begin
                state_d = WAIT_HALF;
            end
        end
    endcase
end

always @(posedge clk) begin
    if (rst) begin
        ctr_q <= 3'b0;
        data_q <= 8'b0;
        sck_q <= 4'b0;
        mosi_q <= 1'b0;
        state_q <= IDLE;
        data_out_q <= 8'b0;
        new_data_q <= 1'b0;
    end else begin
        ctr_q <= ctr_d;
        data_q <= data_d;
        sck_q <= sck_d;
        mosi_q <= mosi_d;
        state_q <= state_d;
        data_out_q <= data_out_d;
        new_data_q <= new_data_d;
    end
end

endmodule
